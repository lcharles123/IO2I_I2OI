module Int_Mul_ALU();

endmodule

module Finished_Store_Buffer();

endmodule

module Issue();

endmodule


module Score_Board();

endmodule

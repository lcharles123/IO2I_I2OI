module Issue_Queue
(
	input clk, rst, stall,
	input [31:0] d_pc, d_sigext,  // Imm
	input [5:0] d_opcode, //adicao de opcode
	input [4:0] d_inst1, d_inst2, d_inst3, 
	
	output reg [31:0] e_pc, e_sigext, // Imm
	output reg [5:0] e_opcode, //adicao de opcode
	output reg [4:0] e_inst1, e_inst2, e_inst3,
	output cheio
);
	reg [5:0] 	pc 	[0:7]; //posicao da instrucao atual
	
	reg [5:0] 	opcode 	[0:7]; //o IQ tera 8 entradas, 6 bits para o opcode
	reg [31:0] 	imm 	[0:7]; // 32 bits para sigext == imm
 
	reg [1:0] 	v 		[0:7]; //se o dest eh valido(todas exceto branch e store)
	reg [4:0] 	dest  	[0:7]; //endDest do banco de regs
	
	reg [1:0] 	v1 		[0:7]; //se fonte0 eh valido
	reg [1:0]	p1 		[0:7];//se fonte0 esta pendente
	reg [5:0]	fonte1 	[0:7];//end fonte0
 
	reg [1:0]	v2 		[0:7];//se fonte1 eh valido
	reg [1:0]	p2 		[0:7];//se fonte1 esta pendente
	reg [5:0] 	fonte2 	[0:7];//end fonte1
	
	reg [1:2] indice_inst_antiga; //guarda o indice da entrada
	reg [1:2] indice_inst_pronta; //guarda o indice da entrada
	reg [1:2] indice_inst_mais_recente; //guarda o indice da entrada
	reg [1:2] contador; //se ==7 , esta cheio	
	
	assign cheio = (contador == 7) ? 1 : 0;
	
//Op: Opcode
//Imm: Imediato
//S: bit especulativo
//V: Válido (Existe no Src e Dest)
//P: Pendente

	always @(posedge clk) 
	begin
      if (!rst) 
		begin
			e_pc       <= 0;
			e_sigext   <= 0;
			e_opcode   <= 0;
			e_inst1    <= 0;
			e_inst2    <= 0;
			e_inst3    <= 0;

			contador				    <= 0;
			indice_inst_antiga   		<= 0; 
			indice_inst_pronta  		<= 0; 
			indice_inst_mais_recente	<= 0;
		end
		else
		begin
			if(!cheio)
			begin
				opcode[indice_inst_mais_recente] = d_opcode;

				imm[indice_inst_mais_recente] = d_sigext;
			
				v[indice_inst_mais_recente] = ~(d_branch || d_memwrite); //se branch ou store -> dest nao valido
				dest[indice_inst_mais_recente] = d_inst3; //endDest do banco de regs

				v1[indice_inst_mais_recente]  = 1; //se fonte1 eh valido
				p1[indice_inst_mais_recente]  = stall;//se fonte1 esta pendente
				fonte1[indice_inst_mais_recente] = d_inst1;//end fonte1
		
				v2[indice_inst_mais_recente]  = 1;//fonte1 eh valido em todos (pois nao tem BEQ por exemplo)
				p2[indice_inst_mais_recente]  = stall;//se fonte2 esta pendente
				fonte2[indice_inst_mais_recente] = (opcode == 6'b000001) ? d_inst3 : d_inst2;//apenas opcode define fonte2
			
				indice_inst_mais_recente = indice_inst_mais_recente + 1;
				contador = contador + 1;
				if(indice_inst_mais_recente == 8)	indice_inst_mais_recente = 0;
			
			end
		
			//Instrucao Pronta = (!VSrc0 || !PSrc0) && (!VSrc1 || !PSrc1) && Sem Hazard Estrutural

			if( (!v1[indice_inst_antiga] || !p1[indice_inst_antiga]) && (!v2[indice_inst_antiga] || !p2[indice_inst_antiga]) && !stall))
			begin
				//envia a instrucao para o issue
				//e_pc       <= ?;
				e_sigext   <= imm[indice_inst_antiga];
				e_opcode   <= opcode[indice_inst_antiga];
				e_inst1    <= fonte1[indice_inst_antiga];
				e_inst2    <= fonte2[indice_inst_antiga];
				e_inst3    <= dest[indice_inst_antiga];
			
				//atualiza os indices
				if(indice_inst_antiga == indice_inst_pronta) indice_inst_pronta = indice_inst_pronta + 1;
				
				indice_inst_antiga = indice_inst_antiga + 1;
				
				if(indice_inst_antiga == 8) indice_inst_antiga = 0;
				
				contador = contador - 1;

			end
			else if((!v1[indice_inst_pronta] || !p1[indice_inst_pronta]) && (!v2[indice_inst_pronta] || !p2[indice_inst_pronta]) && !stall))
			begin
				//envia a instrucao para o issue
				//e_pc       <= ?;
				e_sigext   <= imm[indice_inst_pronta];
				e_opcode   <= opcode[indice_inst_pronta];
				e_inst1    <= fonte1[indice_inst_pronta];
				e_inst2    <= fonte2[indice_inst_pronta];
				e_inst3    <= dest[indice_inst_pronta];
			
				//atualiza os indices
				indice_inst_pronta = indice_inst_pronta + 1;
				
				if(indice_inst_pronta == 8) indice_inst_pronta = 0;

				contador = contador - 1;					
			end
			//else
			//begin
		
			//end	
		end
endmodule

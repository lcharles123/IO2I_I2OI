module Reorder_Buffer();

endmodule

module Phisical_Register_file();

endmodule

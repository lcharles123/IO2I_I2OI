module Commit();

endmodule
